(* This module contains the boolean expression evaluation code
   for KodeLlama2 *)

Require Export Ident.

Module Bexp.

End Bexp.

Export Bexp.

